package yapp_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    typedef uvm_config_db#(virtual yapp_if) yapp_vif_config;

    `include "./sv/yapp_packet.sv"
    `include "./sv/yapp_tx_monitor.sv"
    `include "./sv/yapp_tx_sequencer.sv"
    `include "./sv/yapp_tx_seqs.sv"
    `include "./sv/yapp_tx_driver.sv"
    `include "./sv/yapp_tx_agent.sv"
    `include "./sv/yapp_tx_env.sv"

endpackage: yapp_pkg